module sj (/*AUTOARG*/);
   output sj__zzdl__sig0;
   output sj__zzdl__sig1;
   output sj__zzdl__sig2;
endmodule
