module sub_b (/*AUTOARG*/);
   output sub_b__top__s1;
   input  sub_a__sub_b__s1;
   input  ssub_b__sub_b__s1_temp;
   
   /*AUTOREG*/
   /*AUTOWIRE*/

endmodule
