`ifndef CLOCK_IF__SV 
`define CLOCK_IF__SV 
interface clock_if();
   logic clk;     // clock 
endinterface
`endif 
