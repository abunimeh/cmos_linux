module ssub_a (/*AUTOARG*/);
   output ssub_a__ssub_b__s1;
   input  top__ssub_a__s2;
   
   /*AUTOREG*/
   /*AUTOWIRE*/
   
endmodule // ssub1
