module top (/*AUTOARG*/);

   /*AUTOREG*/
   /*AUTOWIRE*/

   /* sj AUTO_TEMPLATE (
    .sj__zzdl__\(.*\) (sj@__zzdl__\1),
    );*/
   
   sj #(/*AUTOINSTPARAM*/) sj0 (
                                // .a (b);
                                /*AUTOINST*/);
   sj #(/*AUTOINSTPARAM*/)sj2 (/*AUTOINST*/);
   zzdl #(/*AUTOINSTPARAM*/) u_zzdl(/*AUTOINST*/);

endmodule // top
// Local Variables:
// verilog-library-directories:(".")
// End:
