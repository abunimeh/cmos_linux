Count(1)
 u_core.ao486_inst.pipeline_inst.read_inst.read_commands_inst.rd_glob_descriptor_value[31:0]
 u_core.ao486_inst.pipeline_inst.read_inst.rd_glob_descriptor_value[31:0]

Count(2)
 u_core.ao486_inst.pipeline_inst.read_inst.read_commands_inst.rd_glob_descriptor_value[63:32]
 u_core.ao486_inst.pipeline_inst.read_inst.rd_glob_descriptor_value[63:32]

Count(3)
 u_core.ao486_inst.pipeline_inst.read_inst.read_commands_inst.rd_glob_descriptor_2_value[31:0]
 u_core.ao486_inst.pipeline_inst.read_inst.rd_glob_descriptor_2_value[31:0]

Count(4)
 u_core.ao486_inst.pipeline_inst.read_inst.read_commands_inst.rd_glob_descriptor_2_value[63:32]
 u_core.ao486_inst.pipeline_inst.read_inst.rd_glob_descriptor_2_value[63:32]

Count(5)
 u_core.ao486_inst.pipeline_inst.read_inst.read_commands_inst.rd_glob_param_1_value[31:0]
 u_core.ao486_inst.pipeline_inst.read_inst.rd_glob_param_1_value[31:0]

Count(6)
 u_core.ao486_inst.pipeline_inst.read_inst.read_commands_inst.rd_glob_param_2_value[31:0]
 u_core.ao486_inst.pipeline_inst.read_inst.rd_glob_param_2_value[31:0]

Count(7)
 u_core.ao486_inst.pipeline_inst.read_inst.read_commands_inst.rd_glob_param_3_value[31:0]
 u_core.ao486_inst.pipeline_inst.read_inst.rd_glob_param_3_value[31:0]

Count(8)
 u_core.ao486_inst.pipeline_inst.read_inst.read_commands_inst.rd_glob_param_4_value[31:0]
 u_core.ao486_inst.pipeline_inst.read_inst.rd_glob_param_4_value[31:0]

Count(9)
 u_core.ao486_inst.pipeline_inst.read_inst.read_commands_inst.rd_glob_param_5_value[31:0]
 u_core.ao486_inst.pipeline_inst.read_inst.rd_glob_param_5_value[31:0]

Count(10)
 u_core.ao486_inst.pipeline_inst.read_inst.read_commands_inst.rd_extra_wire[31:0]
 u_core.ao486_inst.pipeline_inst.read_inst.rd_extra_wire[31:0]

Count(11)
 u_core.ao486_inst.pipeline_inst.read_inst.read_effective_address_inst.rd_address_effective[31:0]
 u_core.ao486_inst.pipeline_inst.read_inst.rd_address_effective[31:0]

Count(12)
 u_core.ao486_inst.pipeline_inst.read_inst.read_commands_inst.io_read_address[15:0]
 u_core.ao486_inst.pipeline_inst.read_inst.io_read_address[15:0]

Count(13)
 u_core.ao486_inst.pipeline_inst.read_inst.read_commands_inst.rd_io_allow_fault
 u_core.ao486_inst.pipeline_inst.read_inst.rd_io_allow_fault

Count(14)
 u_core.ao486_inst.pipeline_inst.read_inst.read_commands_inst.rd_ss_esp_from_tss_fault
 u_core.ao486_inst.pipeline_inst.read_inst.rd_ss_esp_from_tss_fault

Count(15)
 u_core.ao486_inst.pipeline_inst.read_inst.read_commands_inst.rd_glob_descriptor_set
 u_core.ao486_inst.pipeline_inst.read_inst.rd_glob_descriptor_set

Count(16)
 u_core.ao486_inst.pipeline_inst.read_inst.read_commands_inst.rd_glob_descriptor_2_set
 u_core.ao486_inst.pipeline_inst.read_inst.rd_glob_descriptor_2_set

Count(17)
 u_core.ao486_inst.pipeline_inst.read_inst.read_commands_inst.rd_glob_param_1_set
 u_core.ao486_inst.pipeline_inst.read_inst.rd_glob_param_1_set

Count(18)
 u_core.ao486_inst.pipeline_inst.read_inst.read_commands_inst.rd_glob_param_2_set
 u_core.ao486_inst.pipeline_inst.read_inst.rd_glob_param_2_set

Count(19)
 u_core.ao486_inst.pipeline_inst.read_inst.read_commands_inst.rd_glob_param_3_set
 u_core.ao486_inst.pipeline_inst.read_inst.rd_glob_param_3_set

Count(20)
 u_core.ao486_inst.pipeline_inst.read_inst.read_commands_inst.rd_glob_param_4_set
 u_core.ao486_inst.pipeline_inst.read_inst.rd_glob_param_4_set

Count(21)
 u_core.ao486_inst.pipeline_inst.read_inst.read_commands_inst.rd_glob_param_5_set
 u_core.ao486_inst.pipeline_inst.read_inst.rd_glob_param_5_set

Count(22)
 u_core.ao486_inst.pipeline_inst.read_inst.read_commands_inst.rd_dst_is_reg
 u_core.ao486_inst.pipeline_inst.read_inst.rd_dst_is_reg

Count(23)
 u_core.ao486_inst.pipeline_inst.read_inst.read_commands_inst.rd_dst_is_rm
 u_core.ao486_inst.pipeline_inst.read_inst.rd_dst_is_rm

Count(24)
 u_core.ao486_inst.pipeline_inst.read_inst.read_commands_inst.rd_dst_is_memory
 u_core.ao486_inst.pipeline_inst.read_inst.rd_dst_is_memory

Count(25)
 u_core.ao486_inst.pipeline_inst.read_inst.read_commands_inst.rd_dst_is_eax
 u_core.ao486_inst.pipeline_inst.read_inst.rd_dst_is_eax

Count(26)
 u_core.ao486_inst.pipeline_inst.read_inst.read_commands_inst.rd_dst_is_edx_eax
 u_core.ao486_inst.pipeline_inst.read_inst.rd_dst_is_edx_eax

Count(27)
 u_core.ao486_inst.pipeline_inst.read_inst.read_commands_inst.rd_dst_is_implicit_reg
 u_core.ao486_inst.pipeline_inst.read_inst.rd_dst_is_implicit_reg

Count(28)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_glob_descriptor_value[31:0]
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_glob_descriptor_value[31:0]

Count(29)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_glob_descriptor_value[63:32]
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_glob_descriptor_value[63:32]

Count(30)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_glob_descriptor_2_value[31:0]
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_glob_descriptor_2_value[31:0]

Count(31)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_glob_descriptor_2_value[63:32]
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_glob_descriptor_2_value[63:32]

Count(32)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.tlbcheck_address[31:0]
 u_core.ao486_inst.pipeline_inst.execute_inst.tlbcheck_address[31:0]

Count(33)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.tlbflushsingle_address[31:0]
 u_core.ao486_inst.pipeline_inst.execute_inst.tlbflushsingle_address[31:0]

Count(34)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_glob_param_1_value[31:0]
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_glob_param_1_value[31:0]

Count(35)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_glob_param_2_value[31:0]
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_glob_param_2_value[31:0]

Count(36)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_glob_param_3_value[31:0]
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_glob_param_3_value[31:0]

Count(37)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.task_eip[31:0]
 u_core.ao486_inst.pipeline_inst.execute_inst.task_eip[31:0]

Count(38)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_buffer[31:0]
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_buffer[31:0]

Count(39)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_result[31:0]
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_result[31:0]

Count(40)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_result2[31:0]
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_result2[31:0]

Count(41)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_result_push[31:0]
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_result_push[31:0]

Count(42)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_offset_inst.exe_stack_offset[31:0]
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_stack_offset[31:0]

Count(43)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_buffer_shifted[31:0]
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_buffer_shifted[31:0]

Count(44)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_buffer_shifted[63:32]
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_buffer_shifted[63:32]

Count(45)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_buffer_shifted[95:64]
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_buffer_shifted[95:64]

Count(46)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_buffer_shifted[127:96]
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_buffer_shifted[127:96]

Count(47)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_buffer_shifted[159:128]
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_buffer_shifted[159:128]

Count(48)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_buffer_shifted[191:160]
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_buffer_shifted[191:160]

Count(49)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_buffer_shifted[223:192]
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_buffer_shifted[223:192]

Count(50)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_buffer_shifted[255:224]
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_buffer_shifted[255:224]

Count(51)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_buffer_shifted[287:256]
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_buffer_shifted[287:256]

Count(52)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_buffer_shifted[319:288]
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_buffer_shifted[319:288]

Count(53)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_buffer_shifted[351:320]
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_buffer_shifted[351:320]

Count(54)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_buffer_shifted[383:352]
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_buffer_shifted[383:352]

Count(55)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_buffer_shifted[415:384]
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_buffer_shifted[415:384]

Count(56)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_buffer_shifted[447:416]
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_buffer_shifted[447:416]

Count(57)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_buffer_shifted[463:448]
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_buffer_shifted[463:448]

Count(58)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_result_signals[4:0]
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_result_signals[4:0]

Count(59)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_arith_index[3:0]
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_arith_index[3:0]

Count(60)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.tlbcheck_do
 u_core.ao486_inst.pipeline_inst.execute_inst.tlbcheck_do

Count(61)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.tlbcheck_rw
 u_core.ao486_inst.pipeline_inst.execute_inst.tlbcheck_rw

Count(62)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.tlbflushsingle_do
 u_core.ao486_inst.pipeline_inst.execute_inst.tlbflushsingle_do

Count(63)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.invdcode_do
 u_core.ao486_inst.pipeline_inst.execute_inst.invdcode_do

Count(64)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.invddata_do
 u_core.ao486_inst.pipeline_inst.execute_inst.invddata_do

Count(65)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.wbinvddata_do
 u_core.ao486_inst.pipeline_inst.execute_inst.wbinvddata_do

Count(66)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_glob_descriptor_set
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_glob_descriptor_set

Count(67)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_glob_descriptor_2_set
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_glob_descriptor_2_set

Count(68)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_glob_param_1_set
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_glob_param_1_set

Count(69)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_glob_param_2_set
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_glob_param_2_set

Count(70)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_glob_param_3_set
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_glob_param_3_set

Count(71)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.dr6_bd_set
 u_core.ao486_inst.pipeline_inst.execute_inst.dr6_bd_set

Count(72)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_bound_fault
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_bound_fault

Count(73)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_trigger_gp_fault
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_trigger_gp_fault

Count(74)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_trigger_ts_fault
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_trigger_ts_fault

Count(75)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_trigger_ss_fault
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_trigger_ss_fault

Count(76)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_trigger_np_fault
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_trigger_np_fault

Count(77)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_trigger_pf_fault
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_trigger_pf_fault

Count(78)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_trigger_db_fault
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_trigger_db_fault

Count(79)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_trigger_nm_fault
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_trigger_nm_fault

Count(80)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_load_seg_gp_fault
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_load_seg_gp_fault

Count(81)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_load_seg_ss_fault
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_load_seg_ss_fault

Count(82)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_load_seg_np_fault
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_load_seg_np_fault

Count(83)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_arith_sub_carry
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_arith_sub_carry

Count(84)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_arith_add_carry
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_arith_add_carry

Count(85)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_arith_adc_carry
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_arith_adc_carry

Count(86)
 u_core.ao486_inst.pipeline_inst.execute_inst.execute_commands_inst.exe_arith_sbb_carry
 u_core.ao486_inst.pipeline_inst.execute_inst.exe_arith_sbb_carry

Count(87)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.es_cache[31:0]
 u_core.ao486_inst.pipeline_inst.write_inst.es_cache[31:0]

Count(88)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.es_cache[63:32]
 u_core.ao486_inst.pipeline_inst.write_inst.es_cache[63:32]

Count(89)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.ds_cache[31:0]
 u_core.ao486_inst.pipeline_inst.write_inst.ds_cache[31:0]

Count(90)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.ds_cache[63:32]
 u_core.ao486_inst.pipeline_inst.write_inst.ds_cache[63:32]

Count(91)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.ss_cache[31:0]
 u_core.ao486_inst.pipeline_inst.write_inst.ss_cache[31:0]

Count(92)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.ss_cache[63:32]
 u_core.ao486_inst.pipeline_inst.write_inst.ss_cache[63:32]

Count(93)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.fs_cache[31:0]
 u_core.ao486_inst.pipeline_inst.write_inst.fs_cache[31:0]

Count(94)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.fs_cache[63:32]
 u_core.ao486_inst.pipeline_inst.write_inst.fs_cache[63:32]

Count(95)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.gs_cache[31:0]
 u_core.ao486_inst.pipeline_inst.write_inst.gs_cache[31:0]

Count(96)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.gs_cache[63:32]
 u_core.ao486_inst.pipeline_inst.write_inst.gs_cache[63:32]

Count(97)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.cs_cache[31:0]
 u_core.ao486_inst.pipeline_inst.write_inst.cs_cache[31:0]

Count(98)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.cs_cache[63:32]
 u_core.ao486_inst.pipeline_inst.write_inst.cs_cache[63:32]

Count(99)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.ldtr_cache[31:0]
 u_core.ao486_inst.pipeline_inst.write_inst.ldtr_cache[31:0]

Count(100)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.ldtr_cache[63:32]
 u_core.ao486_inst.pipeline_inst.write_inst.ldtr_cache[63:32]

Count(101)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.tr_cache[31:0]
 u_core.ao486_inst.pipeline_inst.write_inst.tr_cache[31:0]

Count(102)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.tr_cache[63:32]
 u_core.ao486_inst.pipeline_inst.write_inst.tr_cache[63:32]

Count(103)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.gdtr_base[31:0]
 u_core.ao486_inst.pipeline_inst.write_inst.gdtr_base[31:0]

Count(104)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.idtr_base[31:0]
 u_core.ao486_inst.pipeline_inst.write_inst.idtr_base[31:0]

Count(105)
 u_core.ao486_inst.pipeline_inst.write_inst.write_commands_inst.wr_glob_param_1_value[31:0]
 u_core.ao486_inst.pipeline_inst.write_inst.wr_glob_param_1_value[31:0]

Count(106)
 u_core.ao486_inst.pipeline_inst.write_inst.write_commands_inst.wr_glob_param_3_value[31:0]
 u_core.ao486_inst.pipeline_inst.write_inst.wr_glob_param_3_value[31:0]

Count(107)
 u_core.ao486_inst.pipeline_inst.write_inst.write_commands_inst.wr_glob_param_4_value[31:0]
 u_core.ao486_inst.pipeline_inst.write_inst.wr_glob_param_4_value[31:0]

Count(108)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.eax[31:0]
 u_core.ao486_inst.pipeline_inst.write_inst.eax[31:0]

Count(109)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.ebx[31:0]
 u_core.ao486_inst.pipeline_inst.write_inst.ebx[31:0]

Count(110)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.ecx[31:0]
 u_core.ao486_inst.pipeline_inst.write_inst.ecx[31:0]

Count(111)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.edx[31:0]
 u_core.ao486_inst.pipeline_inst.write_inst.edx[31:0]

Count(112)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.esi[31:0]
 u_core.ao486_inst.pipeline_inst.write_inst.esi[31:0]

Count(113)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.edi[31:0]
 u_core.ao486_inst.pipeline_inst.write_inst.edi[31:0]

Count(114)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.ebp[31:0]
 u_core.ao486_inst.pipeline_inst.write_inst.ebp[31:0]

Count(115)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.esp[31:0]
 u_core.ao486_inst.pipeline_inst.write_inst.esp[31:0]

Count(116)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.cr2[31:0]
 u_core.ao486_inst.pipeline_inst.write_inst.cr2[31:0]

Count(117)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.cr3[31:0]
 u_core.ao486_inst.pipeline_inst.write_inst.cr3[31:0]

Count(118)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.dr0[31:0]
 u_core.ao486_inst.pipeline_inst.write_inst.dr0[31:0]

Count(119)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.dr1[31:0]
 u_core.ao486_inst.pipeline_inst.write_inst.dr1[31:0]

Count(120)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.dr2[31:0]
 u_core.ao486_inst.pipeline_inst.write_inst.dr2[31:0]

Count(121)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.dr3[31:0]
 u_core.ao486_inst.pipeline_inst.write_inst.dr3[31:0]

Count(122)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.dr7[31:0]
 u_core.ao486_inst.pipeline_inst.write_inst.dr7[31:0]

Count(123)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.gdtr_limit[15:0]
 u_core.ao486_inst.pipeline_inst.write_inst.gdtr_limit[15:0]

Count(124)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.idtr_limit[15:0]
 u_core.ao486_inst.pipeline_inst.write_inst.idtr_limit[15:0]

Count(125)
 u_core.ao486_inst.pipeline_inst.write_inst.write_commands_inst.wr_error_code[15:0]
 u_core.ao486_inst.pipeline_inst.write_inst.wr_error_code[15:0]

Count(126)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.es[15:0]
 u_core.ao486_inst.pipeline_inst.write_inst.es[15:0]

Count(127)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.ds[15:0]
 u_core.ao486_inst.pipeline_inst.write_inst.ds[15:0]

Count(128)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.ss[15:0]
 u_core.ao486_inst.pipeline_inst.write_inst.ss[15:0]

Count(129)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.fs[15:0]
 u_core.ao486_inst.pipeline_inst.write_inst.fs[15:0]

Count(130)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.gs[15:0]
 u_core.ao486_inst.pipeline_inst.write_inst.gs[15:0]

Count(131)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.cs[15:0]
 u_core.ao486_inst.pipeline_inst.write_inst.cs[15:0]

Count(132)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.ldtr[15:0]
 u_core.ao486_inst.pipeline_inst.write_inst.ldtr[15:0]

Count(133)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.tr[15:0]
 u_core.ao486_inst.pipeline_inst.write_inst.tr[15:0]

Count(134)
 u_core.ao486_inst.pipeline_inst.write_inst.write_commands_inst.wr_int_vector[7:0]
 u_core.ao486_inst.pipeline_inst.write_inst.wr_int_vector[7:0]

Count(135)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.dr6_breakpoints[3:0]
 u_core.ao486_inst.pipeline_inst.write_inst.dr6_breakpoints[3:0]

Count(136)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.debug_len0[2:0]
 u_core.ao486_inst.pipeline_inst.write_inst.debug_len0[2:0]

Count(137)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.debug_len2[2:0]
 u_core.ao486_inst.pipeline_inst.write_inst.debug_len2[2:0]

Count(138)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.debug_len3[2:0]
 u_core.ao486_inst.pipeline_inst.write_inst.debug_len3[2:0]

Count(139)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.cpl[1:0]
 u_core.ao486_inst.pipeline_inst.write_inst.cpl[1:0]

Count(140)
 u_core.ao486_inst.pipeline_inst.write_inst.write_commands_inst.wr_task_rpl[1:0]
 u_core.ao486_inst.pipeline_inst.write_inst.wr_task_rpl[1:0]

Count(141)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.iopl[1:0]
 u_core.ao486_inst.pipeline_inst.write_inst.iopl[1:0]

Count(142)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.real_mode
 u_core.ao486_inst.pipeline_inst.write_inst.real_mode

Count(143)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.v8086_mode
 u_core.ao486_inst.pipeline_inst.write_inst.v8086_mode

Count(144)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.protected_mode
 u_core.ao486_inst.pipeline_inst.write_inst.protected_mode

Count(145)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.io_allow_check_needed
 u_core.ao486_inst.pipeline_inst.write_inst.io_allow_check_needed

Count(146)
 u_core.ao486_inst.pipeline_inst.write_inst.write_commands_inst.wr_int
 u_core.ao486_inst.pipeline_inst.write_inst.wr_int

Count(147)
 u_core.ao486_inst.pipeline_inst.write_inst.write_commands_inst.wr_int_soft_int
 u_core.ao486_inst.pipeline_inst.write_inst.wr_int_soft_int

Count(148)
 u_core.ao486_inst.pipeline_inst.write_inst.write_commands_inst.wr_int_soft_int_ib
 u_core.ao486_inst.pipeline_inst.write_inst.wr_int_soft_int_ib

Count(149)
 u_core.ao486_inst.pipeline_inst.write_inst.write_commands_inst.wr_exception_external_set
 u_core.ao486_inst.pipeline_inst.write_inst.wr_exception_external_set

Count(150)
 u_core.ao486_inst.pipeline_inst.write_inst.write_commands_inst.wr_exception_finished
 u_core.ao486_inst.pipeline_inst.write_inst.wr_exception_finished

Count(151)
 u_core.ao486_inst.pipeline_inst.write_inst.write_stack_inst.wr_new_push_ss_fault
 u_core.ao486_inst.pipeline_inst.write_inst.wr_new_push_ss_fault

Count(152)
 u_core.ao486_inst.pipeline_inst.write_inst.write_string_inst.wr_string_es_fault
 u_core.ao486_inst.pipeline_inst.write_inst.wr_string_es_fault

Count(153)
 u_core.ao486_inst.pipeline_inst.write_inst.write_stack_inst.wr_push_ss_fault
 u_core.ao486_inst.pipeline_inst.write_inst.wr_push_ss_fault

Count(154)
 u_core.ao486_inst.pipeline_inst.write_inst.write_commands_inst.wr_req_reset_pr
 u_core.ao486_inst.pipeline_inst.write_inst.wr_req_reset_pr

Count(155)
 u_core.ao486_inst.pipeline_inst.write_inst.write_commands_inst.wr_req_reset_dec
 u_core.ao486_inst.pipeline_inst.write_inst.wr_req_reset_dec

Count(156)
 u_core.ao486_inst.pipeline_inst.write_inst.write_commands_inst.wr_req_reset_micro
 u_core.ao486_inst.pipeline_inst.write_inst.wr_req_reset_micro

Count(157)
 u_core.ao486_inst.pipeline_inst.write_inst.write_commands_inst.wr_req_reset_rd
 u_core.ao486_inst.pipeline_inst.write_inst.wr_req_reset_rd

Count(158)
 u_core.ao486_inst.pipeline_inst.write_inst.write_commands_inst.wr_req_reset_exe
 u_core.ao486_inst.pipeline_inst.write_inst.wr_req_reset_exe

Count(159)
 u_core.ao486_inst.pipeline_inst.write_inst.write_commands_inst.tlbflushall_do
 u_core.ao486_inst.pipeline_inst.write_inst.tlbflushall_do

Count(160)
 u_core.ao486_inst.pipeline_inst.write_inst.write_commands_inst.wr_glob_param_1_set
 u_core.ao486_inst.pipeline_inst.write_inst.wr_glob_param_1_set

Count(161)
 u_core.ao486_inst.pipeline_inst.write_inst.write_commands_inst.wr_glob_param_3_set
 u_core.ao486_inst.pipeline_inst.write_inst.wr_glob_param_3_set

Count(162)
 u_core.ao486_inst.pipeline_inst.write_inst.write_commands_inst.wr_glob_param_4_set
 u_core.ao486_inst.pipeline_inst.write_inst.wr_glob_param_4_set

Count(163)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.cr0_pe
 u_core.ao486_inst.pipeline_inst.write_inst.cr0_pe

Count(164)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.cr0_mp
 u_core.ao486_inst.pipeline_inst.write_inst.cr0_mp

Count(165)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.cr0_em
 u_core.ao486_inst.pipeline_inst.write_inst.cr0_em

Count(166)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.cr0_ts
 u_core.ao486_inst.pipeline_inst.write_inst.cr0_ts

Count(167)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.cr0_ne
 u_core.ao486_inst.pipeline_inst.write_inst.cr0_ne

Count(168)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.cr0_wp
 u_core.ao486_inst.pipeline_inst.write_inst.cr0_wp

Count(169)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.cr0_am
 u_core.ao486_inst.pipeline_inst.write_inst.cr0_am

Count(170)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.cr0_nw
 u_core.ao486_inst.pipeline_inst.write_inst.cr0_nw

Count(171)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.cr0_cd
 u_core.ao486_inst.pipeline_inst.write_inst.cr0_cd

Count(172)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.cr0_pg
 u_core.ao486_inst.pipeline_inst.write_inst.cr0_pg

Count(173)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.cflag
 u_core.ao486_inst.pipeline_inst.write_inst.cflag

Count(174)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.pflag
 u_core.ao486_inst.pipeline_inst.write_inst.pflag

Count(175)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.aflag
 u_core.ao486_inst.pipeline_inst.write_inst.aflag

Count(176)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.zflag
 u_core.ao486_inst.pipeline_inst.write_inst.zflag

Count(177)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.sflag
 u_core.ao486_inst.pipeline_inst.write_inst.sflag

Count(178)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.oflag
 u_core.ao486_inst.pipeline_inst.write_inst.oflag

Count(179)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.tflag
 u_core.ao486_inst.pipeline_inst.write_inst.tflag

Count(180)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.iflag
 u_core.ao486_inst.pipeline_inst.write_inst.iflag

Count(181)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.dflag
 u_core.ao486_inst.pipeline_inst.write_inst.dflag

Count(182)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.ntflag
 u_core.ao486_inst.pipeline_inst.write_inst.ntflag

Count(183)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.rflag
 u_core.ao486_inst.pipeline_inst.write_inst.rflag

Count(184)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.vmflag
 u_core.ao486_inst.pipeline_inst.write_inst.vmflag

Count(185)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.acflag
 u_core.ao486_inst.pipeline_inst.write_inst.acflag

Count(186)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.idflag
 u_core.ao486_inst.pipeline_inst.write_inst.idflag

Count(187)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.dr6_b12
 u_core.ao486_inst.pipeline_inst.write_inst.dr6_b12

Count(188)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.dr6_bd
 u_core.ao486_inst.pipeline_inst.write_inst.dr6_bd

Count(189)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.dr6_bs
 u_core.ao486_inst.pipeline_inst.write_inst.dr6_bs

Count(190)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.dr6_bt
 u_core.ao486_inst.pipeline_inst.write_inst.dr6_bt

Count(191)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.es_cache_valid
 u_core.ao486_inst.pipeline_inst.write_inst.es_cache_valid

Count(192)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.ds_cache_valid
 u_core.ao486_inst.pipeline_inst.write_inst.ds_cache_valid

Count(193)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.ss_cache_valid
 u_core.ao486_inst.pipeline_inst.write_inst.ss_cache_valid

Count(194)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.fs_cache_valid
 u_core.ao486_inst.pipeline_inst.write_inst.fs_cache_valid

Count(195)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.gs_cache_valid
 u_core.ao486_inst.pipeline_inst.write_inst.gs_cache_valid

Count(196)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.cs_cache_valid
 u_core.ao486_inst.pipeline_inst.write_inst.cs_cache_valid

Count(197)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.ldtr_cache_valid
 u_core.ao486_inst.pipeline_inst.write_inst.ldtr_cache_valid

Count(198)
 u_core.ao486_inst.pipeline_inst.write_inst.write_register_inst.tr_cache_valid
 u_core.ao486_inst.pipeline_inst.write_inst.tr_cache_valid

Count(199)
 u_core.ao486_inst.memory_inst.avalon_mem_inst.avm_address[31:0]
 u_core.ao486_inst.avm_address[31:0]

Count(200)
 u_core.ao486_inst.memory_inst.avalon_mem_inst.avm_writedata[31:0]
 u_core.ao486_inst.avm_writedata[31:0]

Count(201)
 u_core.ao486_inst.avalon_io_inst.avalon_io_writedata[31:0]
 u_core.ao486_inst.avalon_io_writedata[31:0]

Count(202)
 u_core.ao486_inst.avalon_io_inst.avalon_io_address[15:0]
 u_core.ao486_inst.avalon_io_address[15:0]

Count(203)
 u_core.ao486_inst.memory_inst.avalon_mem_inst.avm_byteenable[3:0]
 u_core.ao486_inst.avm_byteenable[3:0]

Count(204)
 u_core.ao486_inst.avalon_io_inst.avalon_io_byteenable[3:0]
 u_core.ao486_inst.avalon_io_byteenable[3:0]

Count(205)
 u_core.ao486_inst.memory_inst.avalon_mem_inst.avm_burstcount[2:0]
 u_core.ao486_inst.avm_burstcount[2:0]

Count(206)
 u_core.ao486_inst.exception_inst.interrupt_done
 u_core.ao486_inst.interrupt_done

Count(207)
 u_core.ao486_inst.memory_inst.avalon_mem_inst.avm_write
 u_core.ao486_inst.avm_write

Count(208)
 u_core.ao486_inst.memory_inst.avalon_mem_inst.avm_read
 u_core.ao486_inst.avm_read

Count(209)
 u_core.ao486_inst.avalon_io_inst.avalon_io_read
 u_core.ao486_inst.avalon_io_read

Count(210)
 u_core.ao486_inst.avalon_io_inst.avalon_io_write
 u_core.ao486_inst.avalon_io_write

The total Count is 210!!!
