module zzdl (/*AUTOARG*/);
   input sj0__zzdl__sig0;
   input sj0__zzdl__sig1;
   input sj0__zzdl__sig2;
   input sj2__zzdl__sig0;
   input sj2__zzdl__sig1;
   input sj2__zzdl__sig2;
endmodule // zzdl
