module ssub_b (/*AUTOARG*/);
   output ssub_b__sub_b__s1;
   input  top__ssub_b__s3;
   input  ssub_a__ssub_b__s1;
   
   /*AUTOREG*/
   /*AUTOWIRE*/
   
endmodule // ssub1
